interface inter;
  
  logic clk;
  logic rd, wr;
  logic full, empty;
  logic [7:0] din;
  logic [7:0] dout;
  logic rst;
  
endinterface
