interface inter(input logic clk);//clock is generating and comming from (testbench.sv) top module so it is input for interface
  //interface has all dut signals
  //Declare with logic type
  //logic clk;
  
  logic rst;
  logic d;
  logic q;
  
endinterface
